package udp_master_pkg;
    
    typedef enum {ARP, Eth2AXI, RAW} type_pkt_t;

endpackage