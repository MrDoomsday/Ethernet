package pkg_decoder;
    // интерфейсы для подключения к портам модуля
    `include "axis_sink.sv"
    `include "axis_source.sv"

    `include "packet.sv"

endpackage