class agent_axis;

    generator_slave gen;
    driver_axis drv;
    monitor_axis mon;
    monitor_mac mon_mac;


    function new();
        gen = new();
        drv = new();
        mon = new();
        mon_mac = new();
    endfunction

    virtual task run();
        fork
            gen.run();
            drv.run();
            mon.run();
            mon_mac.run();
        join
    endtask

endclass


class agent_axim;

    driver_axim drv;
    monitor_axis mon;


    function new();
        drv = new();
        mon = new();
    endfunction

    virtual task run();
        fork
            drv.run();
            mon.run();
        join
    endtask

endclass